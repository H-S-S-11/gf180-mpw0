module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vdd,
    vss,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vdd;
 input vss;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire net114;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net115;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net116;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net85;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net86;
 wire net103;
 wire net104;
 wire net105;
 wire net87;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net21;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net22;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net23;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net24;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net25;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net26;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire \mod.dice0.DiceValue[0] ;
 wire \mod.dice0.DiceValue[1] ;
 wire \mod.dice0.cont1.enable_reg ;
 wire \mod.dice0.rand1.lfsr[0].D ;
 wire \mod.dice0.rand1.lfsr[0].Q ;
 wire \mod.dice0.rand1.lfsr[10].D ;
 wire \mod.dice0.rand1.lfsr[10].Q ;
 wire \mod.dice0.rand1.lfsr[1].D ;
 wire \mod.dice0.rand1.lfsr[2].D ;
 wire \mod.dice0.rand1.lfsr[2].nQ ;
 wire \mod.dice0.rand1.lfsr[3].D ;
 wire \mod.dice0.rand1.lfsr[4].D ;
 wire \mod.dice0.rand1.lfsr[5].D ;
 wire \mod.dice0.rand1.lfsr[6].D ;
 wire \mod.dice0.rand1.lfsr[7].D ;
 wire \mod.dice0.rand1.lfsr[8].D ;
 wire \mod.pdm_core.accumulator[0] ;
 wire \mod.pdm_core.accumulator[1] ;
 wire \mod.pdm_core.accumulator[2] ;
 wire \mod.pdm_core.accumulator[3] ;
 wire \mod.pdm_core.accumulator[4] ;
 wire \mod.pdm_core.input_reg[0] ;
 wire \mod.pdm_core.input_reg[1] ;
 wire \mod.pdm_core.input_reg[2] ;
 wire \mod.pdm_core.input_reg[3] ;
 wire \mod.pdm_core.input_reg[4] ;
 wire \mod.pdm_core.sum[0] ;
 wire \mod.pdm_core.sum[1] ;
 wire \mod.pdm_core.sum[2] ;
 wire \mod.pdm_core.sum[3] ;
 wire \mod.pdm_core.sum[4] ;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net157;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net158;
 wire net186;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;

 gf180mcu_fd_sc_mcu7t5v0__buf_2 _076_ (.I(net1),
    .Z(_047_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _077_ (.I0(\mod.pdm_core.input_reg[4] ),
    .I1(net6),
    .S(_047_),
    .Z(_048_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _078_ (.I(_048_),
    .Z(_016_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _079_ (.I0(\mod.pdm_core.input_reg[3] ),
    .I1(net5),
    .S(_047_),
    .Z(_049_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _080_ (.I(_049_),
    .Z(_015_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _081_ (.I0(\mod.pdm_core.input_reg[2] ),
    .I1(net4),
    .S(_047_),
    .Z(_050_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _082_ (.I(_050_),
    .Z(_014_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _083_ (.I0(\mod.pdm_core.input_reg[1] ),
    .I1(net3),
    .S(_047_),
    .Z(_051_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _084_ (.I(_051_),
    .Z(_013_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _085_ (.I0(\mod.pdm_core.input_reg[0] ),
    .I1(net2),
    .S(net1),
    .Z(_052_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _086_ (.I(_052_),
    .Z(_012_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _087_ (.I(\mod.dice0.cont1.enable_reg ),
    .ZN(_053_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _088_ (.I(_053_),
    .Z(_000_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _089_ (.I(net17),
    .Z(_054_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _090_ (.I(_054_),
    .Z(_055_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _091_ (.I(\mod.dice0.DiceValue[1] ),
    .Z(_056_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _092_ (.A1(_055_),
    .A2(_056_),
    .Z(_057_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _093_ (.I(_057_),
    .Z(net19),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _094_ (.A1(_055_),
    .A2(_056_),
    .Z(_058_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _095_ (.I(_058_),
    .Z(net18),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _096_ (.I(\mod.dice0.DiceValue[0] ),
    .Z(_059_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _097_ (.I(_059_),
    .ZN(_060_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _098_ (.A1(_060_),
    .A2(net18),
    .ZN(net16),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _099_ (.I(\mod.dice0.rand1.lfsr[2].D ),
    .ZN(_001_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _100_ (.A1(\mod.pdm_core.input_reg[4] ),
    .A2(\mod.pdm_core.accumulator[4] ),
    .ZN(_061_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _101_ (.A1(\mod.pdm_core.input_reg[4] ),
    .A2(\mod.pdm_core.accumulator[4] ),
    .Z(_062_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _102_ (.A1(\mod.pdm_core.input_reg[3] ),
    .A2(\mod.pdm_core.accumulator[3] ),
    .ZN(_063_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _103_ (.A1(\mod.pdm_core.input_reg[2] ),
    .A2(\mod.pdm_core.accumulator[2] ),
    .ZN(_064_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _104_ (.A1(\mod.pdm_core.input_reg[0] ),
    .A2(\mod.pdm_core.accumulator[0] ),
    .Z(_065_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _105_ (.A1(\mod.pdm_core.input_reg[1] ),
    .A2(\mod.pdm_core.accumulator[1] ),
    .Z(_066_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _106_ (.A1(\mod.pdm_core.input_reg[1] ),
    .A2(\mod.pdm_core.accumulator[1] ),
    .Z(_067_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _107_ (.A1(\mod.pdm_core.input_reg[2] ),
    .A2(\mod.pdm_core.accumulator[2] ),
    .B1(_065_),
    .B2(_066_),
    .C(_067_),
    .ZN(_068_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _108_ (.A1(\mod.pdm_core.input_reg[3] ),
    .A2(\mod.pdm_core.accumulator[3] ),
    .ZN(_069_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _109_ (.A1(_063_),
    .A2(_064_),
    .A3(_068_),
    .B(_069_),
    .ZN(_070_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _110_ (.A1(_062_),
    .A2(_070_),
    .ZN(_071_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _111_ (.A1(_061_),
    .A2(_071_),
    .ZN(net11),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _112_ (.A1(_061_),
    .A2(_071_),
    .Z(_072_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _113_ (.I(_072_),
    .Z(net12),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _114_ (.I(\mod.dice0.rand1.lfsr[0].Q ),
    .Z(_073_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _115_ (.A1(_073_),
    .A2(\mod.dice0.rand1.lfsr[2].nQ ),
    .Z(_074_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _116_ (.I(_074_),
    .Z(\mod.dice0.rand1.lfsr[10].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _117_ (.A1(\mod.pdm_core.input_reg[0] ),
    .A2(\mod.pdm_core.accumulator[0] ),
    .Z(_075_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _118_ (.I(_075_),
    .Z(\mod.pdm_core.sum[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _119_ (.A1(_065_),
    .A2(_066_),
    .Z(_020_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _120_ (.I(_020_),
    .Z(\mod.pdm_core.sum[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _121_ (.A1(_065_),
    .A2(_066_),
    .B(_067_),
    .ZN(_021_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _122_ (.A1(\mod.pdm_core.input_reg[2] ),
    .A2(\mod.pdm_core.accumulator[2] ),
    .A3(_021_),
    .ZN(_022_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _123_ (.I(_022_),
    .Z(\mod.pdm_core.sum[2] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _124_ (.A1(_064_),
    .A2(_068_),
    .ZN(_023_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _125_ (.A1(\mod.pdm_core.input_reg[3] ),
    .A2(\mod.pdm_core.accumulator[3] ),
    .A3(_023_),
    .Z(_024_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _126_ (.I(_024_),
    .Z(\mod.pdm_core.sum[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _127_ (.A1(_062_),
    .A2(_070_),
    .Z(_025_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _128_ (.I(_025_),
    .Z(\mod.pdm_core.sum[4] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _129_ (.I(net10),
    .Z(_026_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _130_ (.I(_026_),
    .ZN(_002_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _131_ (.I(_026_),
    .ZN(_003_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _132_ (.I(_026_),
    .ZN(_004_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _133_ (.I(_026_),
    .ZN(_005_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _134_ (.I(net10),
    .Z(_027_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _135_ (.I(_027_),
    .ZN(_006_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _136_ (.I(_027_),
    .ZN(_007_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _137_ (.I(_027_),
    .ZN(_008_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _138_ (.I(_027_),
    .ZN(_009_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _139_ (.I(net10),
    .ZN(_010_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _140_ (.I(net10),
    .ZN(_011_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _141_ (.A1(net17),
    .A2(\mod.dice0.DiceValue[1] ),
    .Z(_028_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _142_ (.A1(\mod.dice0.DiceValue[1] ),
    .A2(\mod.dice0.DiceValue[0] ),
    .ZN(_029_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _143_ (.I(\mod.dice0.rand1.lfsr[0].D ),
    .ZN(_030_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _144_ (.A1(_028_),
    .A2(_029_),
    .B(_030_),
    .ZN(_031_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _145_ (.A1(_073_),
    .A2(_031_),
    .B(_053_),
    .ZN(_032_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _146_ (.I(\mod.dice0.rand1.lfsr[0].Q ),
    .ZN(_033_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _147_ (.A1(_030_),
    .A2(_028_),
    .A3(_029_),
    .Z(_034_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _148_ (.I(_056_),
    .ZN(_035_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _149_ (.A1(_054_),
    .A2(_035_),
    .A3(_059_),
    .Z(_036_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _150_ (.A1(_054_),
    .A2(_035_),
    .A3(_059_),
    .ZN(_037_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _151_ (.A1(_031_),
    .A2(_034_),
    .A3(_036_),
    .A4(_037_),
    .ZN(_038_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _152_ (.A1(_035_),
    .A2(_059_),
    .ZN(_039_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _153_ (.A1(_054_),
    .A2(_056_),
    .A3(_060_),
    .ZN(_040_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _154_ (.A1(_055_),
    .A2(_039_),
    .B(_040_),
    .ZN(_041_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _155_ (.A1(\mod.dice0.rand1.lfsr[0].D ),
    .A2(_033_),
    .ZN(_042_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _156_ (.A1(_033_),
    .A2(_038_),
    .B1(_041_),
    .B2(_042_),
    .ZN(_043_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _157_ (.A1(_000_),
    .A2(_060_),
    .B1(_032_),
    .B2(_043_),
    .ZN(_017_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _158_ (.A1(\mod.dice0.rand1.lfsr[0].D ),
    .A2(\mod.dice0.rand1.lfsr[0].Q ),
    .ZN(_044_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _159_ (.A1(_073_),
    .A2(_038_),
    .B1(_041_),
    .B2(_044_),
    .ZN(_045_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _160_ (.A1(_000_),
    .A2(_035_),
    .B1(_032_),
    .B2(_045_),
    .ZN(_018_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _161_ (.A1(_053_),
    .A2(_055_),
    .ZN(_046_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _162_ (.A1(_000_),
    .A2(_073_),
    .B(_046_),
    .ZN(_019_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _163_ (.D(_012_),
    .RN(_002_),
    .CLK(net9),
    .Q(\mod.pdm_core.input_reg[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _164_ (.D(_013_),
    .RN(_003_),
    .CLK(net9),
    .Q(\mod.pdm_core.input_reg[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _165_ (.D(_014_),
    .RN(_004_),
    .CLK(net9),
    .Q(\mod.pdm_core.input_reg[2] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _166_ (.D(_015_),
    .RN(_005_),
    .CLK(net9),
    .Q(\mod.pdm_core.input_reg[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _167_ (.D(_016_),
    .RN(_006_),
    .CLK(net9),
    .Q(\mod.pdm_core.input_reg[4] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _168_ (.D(\mod.dice0.rand1.lfsr[10].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[10].Q ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _169_ (.D(\mod.dice0.rand1.lfsr[10].Q ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[8].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _170_ (.D(\mod.dice0.rand1.lfsr[8].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[7].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _171_ (.D(\mod.dice0.rand1.lfsr[7].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[6].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _172_ (.D(\mod.dice0.rand1.lfsr[6].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[5].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _173_ (.D(\mod.dice0.rand1.lfsr[5].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[4].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _174_ (.D(\mod.dice0.rand1.lfsr[4].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[3].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _175_ (.D(\mod.dice0.rand1.lfsr[3].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[2].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _176_ (.D(\mod.dice0.rand1.lfsr[2].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[1].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _177_ (.D(_001_),
    .SETN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[2].nQ ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _178_ (.D(\mod.dice0.rand1.lfsr[1].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[0].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _179_ (.D(\mod.dice0.rand1.lfsr[0].D ),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.rand1.lfsr[0].Q ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _180_ (.D(_000_),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.cont1.enable_reg ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _181_ (.D(\mod.pdm_core.sum[0] ),
    .RN(_007_),
    .CLK(net9),
    .Q(\mod.pdm_core.accumulator[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _182_ (.D(\mod.pdm_core.sum[1] ),
    .RN(_008_),
    .CLK(net9),
    .Q(\mod.pdm_core.accumulator[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _183_ (.D(\mod.pdm_core.sum[2] ),
    .RN(_009_),
    .CLK(net9),
    .Q(\mod.pdm_core.accumulator[2] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _184_ (.D(\mod.pdm_core.sum[3] ),
    .RN(_010_),
    .CLK(net9),
    .Q(\mod.pdm_core.accumulator[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _185_ (.D(\mod.pdm_core.sum[4] ),
    .RN(_011_),
    .CLK(net9),
    .Q(\mod.pdm_core.accumulator[4] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _186_ (.D(_017_),
    .SETN(net8),
    .CLK(net7),
    .Q(\mod.dice0.DiceValue[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _187_ (.D(_018_),
    .RN(net8),
    .CLK(net7),
    .Q(\mod.dice0.DiceValue[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _188_ (.D(_019_),
    .RN(net8),
    .CLK(net7),
    .Q(net17),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_85 (.ZN(net85),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_86 (.ZN(net86),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_87 (.ZN(net87),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_88 (.ZN(net88),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_89 (.ZN(net89),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_90 (.ZN(net90),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_91 (.ZN(net91),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_92 (.ZN(net92),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_93 (.ZN(net93),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_94 (.ZN(net94),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_95 (.ZN(net95),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_96 (.ZN(net96),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_97 (.ZN(net97),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_98 (.ZN(net98),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_99 (.ZN(net99),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_100 (.ZN(net100),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_101 (.ZN(net101),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_102 (.ZN(net102),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_103 (.ZN(net103),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_104 (.ZN(net104),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_105 (.ZN(net105),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_106 (.ZN(net106),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_107 (.ZN(net107),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_108 (.ZN(net108),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_109 (.ZN(net109),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_110 (.ZN(net110),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_111 (.ZN(net111),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_112 (.ZN(net112),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_113 (.ZN(net113),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_114 (.ZN(net114),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_115 (.ZN(net115),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_116 (.ZN(net116),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_117 (.ZN(net117),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_118 (.ZN(net118),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_119 (.ZN(net119),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_120 (.ZN(net120),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_121 (.ZN(net121),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_122 (.ZN(net122),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_123 (.ZN(net123),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_124 (.ZN(net124),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_125 (.ZN(net125),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_126 (.ZN(net126),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_127 (.ZN(net127),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_128 (.ZN(net128),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_129 (.ZN(net129),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_130 (.ZN(net130),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_131 (.ZN(net131),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_132 (.ZN(net132),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_133 (.ZN(net133),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_134 (.ZN(net134),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_135 (.ZN(net135),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_136 (.ZN(net136),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_137 (.ZN(net137),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_138 (.ZN(net138),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_139 (.ZN(net139),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_140 (.ZN(net140),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_141 (.ZN(net141),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_142 (.ZN(net142),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_143 (.ZN(net143),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_144 (.ZN(net144),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_145 (.ZN(net145),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_146 (.ZN(net146),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_147 (.ZN(net147),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_148 (.ZN(net148),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_149 (.ZN(net149),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_150 (.ZN(net150),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_151 (.ZN(net151),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_152 (.ZN(net152),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_153 (.ZN(net153),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_154 (.ZN(net154),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_155 (.ZN(net155),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_156 (.ZN(net156),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_157 (.ZN(net157),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_158 (.ZN(net158),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_159 (.ZN(net159),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_160 (.ZN(net160),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_161 (.ZN(net161),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_162 (.ZN(net162),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_163 (.ZN(net163),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_164 (.ZN(net164),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_165 (.ZN(net165),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_166 (.ZN(net166),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_167 (.ZN(net167),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_168 (.ZN(net168),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_169 (.ZN(net169),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_170 (.ZN(net170),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_171 (.ZN(net171),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_172 (.ZN(net172),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_173 (.ZN(net173),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_174 (.ZN(net174),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_175 (.ZN(net175),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_176 (.ZN(net176),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_177 (.ZN(net177),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_178 (.ZN(net178),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_179 (.ZN(net179),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_180 (.ZN(net180),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_181 (.ZN(net181),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_182 (.ZN(net182),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_183 (.ZN(net183),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_184 (.ZN(net184),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_185 (.ZN(net185),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_186 (.ZN(net186),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__D (.I(_000_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _356_ (.I(net19),
    .Z(net13),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _357_ (.I(net18),
    .Z(net14),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _358_ (.I(net17),
    .Z(net15),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[10]),
    .Z(net1),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[11]),
    .Z(net2),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[12]),
    .Z(net3),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[13]),
    .Z(net4),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[14]),
    .Z(net5),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[15]),
    .Z(net6),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(io_in[16]),
    .Z(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input8 (.I(io_in[17]),
    .Z(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input9 (.I(io_in[8]),
    .Z(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(io_in[9]),
    .Z(net10),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output11 (.I(net11),
    .Z(io_out[18]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output12 (.I(net12),
    .Z(io_out[19]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output13 (.I(net13),
    .Z(io_out[20]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output14 (.I(net14),
    .Z(io_out[21]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output15 (.I(net15),
    .Z(io_out[22]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output16 (.I(net16),
    .Z(io_out[23]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output17 (.I(net17),
    .Z(io_out[24]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output18 (.I(net18),
    .Z(io_out[25]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output19 (.I(net19),
    .Z(io_out[26]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__A1 (.I(_000_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__A1 (.I(_000_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__A1 (.I(_000_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__RN (.I(_003_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__D (.I(_019_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__I (.I(_025_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__133__I (.I(_026_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__I (.I(_026_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__I (.I(_026_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__130__I (.I(_026_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__I (.I(_027_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__I (.I(_027_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__I (.I(_027_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__I (.I(_027_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__A2 (.I(_028_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__A1 (.I(_028_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__A3 (.I(_029_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__A2 (.I(_029_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__A1 (.I(_030_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__B (.I(_030_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__A1 (.I(_031_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__A2 (.I(_031_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__B1 (.I(_032_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__B1 (.I(_032_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__A1 (.I(_033_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__155__A2 (.I(_033_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__A2 (.I(_035_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__A1 (.I(_035_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__A2 (.I(_035_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__A2 (.I(_035_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__B2 (.I(_042_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__B (.I(_046_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__083__S (.I(_047_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__S (.I(_047_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__S (.I(_047_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__S (.I(_047_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__078__I (.I(_048_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__A1 (.I(_053_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__B (.I(_053_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__I (.I(_053_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__A1 (.I(_054_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__A1 (.I(_054_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__A1 (.I(_054_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__I (.I(_054_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__A2 (.I(_055_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__A1 (.I(_055_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__094__A1 (.I(_055_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__092__A1 (.I(_055_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__A2 (.I(_056_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__I (.I(_056_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__094__A2 (.I(_056_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__092__A2 (.I(_056_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__A2 (.I(_059_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__A3 (.I(_059_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__A3 (.I(_059_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__097__I (.I(_059_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__A2 (.I(_060_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__A3 (.I(_060_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__A1 (.I(_060_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__109__A1 (.I(_063_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__A1 (.I(_064_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__109__A2 (.I(_064_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__A2 (.I(_073_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__A1 (.I(_073_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__A1 (.I(_073_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__115__A1 (.I(_073_),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[14]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[15]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[16]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[17]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[8]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[9]),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A1 (.I(\mod.dice0.DiceValue[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__A2 (.I(\mod.dice0.DiceValue[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__091__I (.I(\mod.dice0.DiceValue[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__D (.I(\mod.dice0.rand1.lfsr[0].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__A1 (.I(\mod.dice0.rand1.lfsr[0].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__155__A1 (.I(\mod.dice0.rand1.lfsr[0].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__I (.I(\mod.dice0.rand1.lfsr[0].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__A2 (.I(\mod.dice0.rand1.lfsr[0].Q ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__I (.I(\mod.dice0.rand1.lfsr[0].Q ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__114__I (.I(\mod.dice0.rand1.lfsr[0].Q ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__D (.I(\mod.dice0.rand1.lfsr[6].D ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__A2 (.I(\mod.pdm_core.accumulator[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__A2 (.I(\mod.pdm_core.accumulator[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__A2 (.I(\mod.pdm_core.accumulator[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A2 (.I(\mod.pdm_core.accumulator[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__A2 (.I(\mod.pdm_core.accumulator[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__A1 (.I(\mod.pdm_core.input_reg[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__A1 (.I(\mod.pdm_core.input_reg[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__085__I0 (.I(\mod.pdm_core.input_reg[0] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__A1 (.I(\mod.pdm_core.input_reg[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__A1 (.I(\mod.pdm_core.input_reg[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__083__I0 (.I(\mod.pdm_core.input_reg[1] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__122__A1 (.I(\mod.pdm_core.input_reg[2] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__A1 (.I(\mod.pdm_core.input_reg[2] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__103__A1 (.I(\mod.pdm_core.input_reg[2] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__I0 (.I(\mod.pdm_core.input_reg[2] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__A1 (.I(\mod.pdm_core.input_reg[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A1 (.I(\mod.pdm_core.input_reg[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__A1 (.I(\mod.pdm_core.input_reg[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__I0 (.I(\mod.pdm_core.input_reg[3] ),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__085__S (.I(net1),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__076__I (.I(net1),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__085__I1 (.I(net2),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__083__I1 (.I(net3),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__I1 (.I(net4),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__I1 (.I(net5),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__I1 (.I(net6),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__CLK (.I(net7),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__SETN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__SETN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__RN (.I(net8),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__CLK (.I(net9),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__I (.I(net10),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__I (.I(net10),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__I (.I(net10),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__I (.I(net10),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__I (.I(net17),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__A1 (.I(net17),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__089__I (.I(net17),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__I (.I(net18),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__A2 (.I(net18),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__I (.I(net19),
    .VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1043 (.VDD(vdd),
    .VSS(vss));
 assign io_oeb[0] = net113;
 assign io_oeb[10] = net123;
 assign io_oeb[11] = net124;
 assign io_oeb[12] = net125;
 assign io_oeb[13] = net126;
 assign io_oeb[14] = net127;
 assign io_oeb[15] = net128;
 assign io_oeb[16] = net129;
 assign io_oeb[17] = net130;
 assign io_oeb[18] = net131;
 assign io_oeb[19] = net132;
 assign io_oeb[1] = net114;
 assign io_oeb[20] = net133;
 assign io_oeb[21] = net134;
 assign io_oeb[22] = net135;
 assign io_oeb[23] = net136;
 assign io_oeb[24] = net137;
 assign io_oeb[25] = net138;
 assign io_oeb[26] = net139;
 assign io_oeb[27] = net140;
 assign io_oeb[28] = net141;
 assign io_oeb[29] = net142;
 assign io_oeb[2] = net115;
 assign io_oeb[30] = net143;
 assign io_oeb[31] = net144;
 assign io_oeb[32] = net145;
 assign io_oeb[33] = net146;
 assign io_oeb[34] = net147;
 assign io_oeb[35] = net148;
 assign io_oeb[36] = net149;
 assign io_oeb[37] = net150;
 assign io_oeb[3] = net116;
 assign io_oeb[4] = net117;
 assign io_oeb[5] = net118;
 assign io_oeb[6] = net119;
 assign io_oeb[7] = net120;
 assign io_oeb[8] = net121;
 assign io_oeb[9] = net122;
 assign io_out[0] = net84;
 assign io_out[10] = net94;
 assign io_out[11] = net95;
 assign io_out[12] = net96;
 assign io_out[13] = net97;
 assign io_out[14] = net98;
 assign io_out[15] = net99;
 assign io_out[16] = net100;
 assign io_out[17] = net101;
 assign io_out[1] = net85;
 assign io_out[27] = net102;
 assign io_out[28] = net103;
 assign io_out[29] = net104;
 assign io_out[2] = net86;
 assign io_out[30] = net105;
 assign io_out[31] = net106;
 assign io_out[32] = net107;
 assign io_out[33] = net108;
 assign io_out[34] = net109;
 assign io_out[35] = net110;
 assign io_out[36] = net111;
 assign io_out[37] = net112;
 assign io_out[3] = net87;
 assign io_out[4] = net88;
 assign io_out[5] = net89;
 assign io_out[6] = net90;
 assign io_out[7] = net91;
 assign io_out[8] = net92;
 assign io_out[9] = net93;
 assign la_data_out[0] = net20;
 assign la_data_out[10] = net30;
 assign la_data_out[11] = net31;
 assign la_data_out[12] = net32;
 assign la_data_out[13] = net33;
 assign la_data_out[14] = net34;
 assign la_data_out[15] = net35;
 assign la_data_out[16] = net36;
 assign la_data_out[17] = net37;
 assign la_data_out[18] = net38;
 assign la_data_out[19] = net39;
 assign la_data_out[1] = net21;
 assign la_data_out[20] = net40;
 assign la_data_out[21] = net41;
 assign la_data_out[22] = net42;
 assign la_data_out[23] = net43;
 assign la_data_out[24] = net44;
 assign la_data_out[25] = net45;
 assign la_data_out[26] = net46;
 assign la_data_out[27] = net47;
 assign la_data_out[28] = net48;
 assign la_data_out[29] = net49;
 assign la_data_out[2] = net22;
 assign la_data_out[30] = net50;
 assign la_data_out[31] = net51;
 assign la_data_out[32] = net52;
 assign la_data_out[33] = net53;
 assign la_data_out[34] = net54;
 assign la_data_out[35] = net55;
 assign la_data_out[36] = net56;
 assign la_data_out[37] = net57;
 assign la_data_out[38] = net58;
 assign la_data_out[39] = net59;
 assign la_data_out[3] = net23;
 assign la_data_out[40] = net60;
 assign la_data_out[41] = net61;
 assign la_data_out[42] = net62;
 assign la_data_out[43] = net63;
 assign la_data_out[44] = net64;
 assign la_data_out[45] = net65;
 assign la_data_out[46] = net66;
 assign la_data_out[47] = net67;
 assign la_data_out[48] = net68;
 assign la_data_out[49] = net69;
 assign la_data_out[4] = net24;
 assign la_data_out[50] = net70;
 assign la_data_out[51] = net71;
 assign la_data_out[52] = net72;
 assign la_data_out[53] = net73;
 assign la_data_out[54] = net74;
 assign la_data_out[55] = net75;
 assign la_data_out[56] = net76;
 assign la_data_out[57] = net77;
 assign la_data_out[58] = net78;
 assign la_data_out[59] = net79;
 assign la_data_out[5] = net25;
 assign la_data_out[60] = net80;
 assign la_data_out[61] = net81;
 assign la_data_out[62] = net82;
 assign la_data_out[63] = net83;
 assign la_data_out[6] = net26;
 assign la_data_out[7] = net27;
 assign la_data_out[8] = net28;
 assign la_data_out[9] = net29;
 assign user_irq[0] = net151;
 assign user_irq[1] = net152;
 assign user_irq[2] = net153;
 assign wbs_ack_o = net154;
 assign wbs_dat_o[0] = net155;
 assign wbs_dat_o[10] = net165;
 assign wbs_dat_o[11] = net166;
 assign wbs_dat_o[12] = net167;
 assign wbs_dat_o[13] = net168;
 assign wbs_dat_o[14] = net169;
 assign wbs_dat_o[15] = net170;
 assign wbs_dat_o[16] = net171;
 assign wbs_dat_o[17] = net172;
 assign wbs_dat_o[18] = net173;
 assign wbs_dat_o[19] = net174;
 assign wbs_dat_o[1] = net156;
 assign wbs_dat_o[20] = net175;
 assign wbs_dat_o[21] = net176;
 assign wbs_dat_o[22] = net177;
 assign wbs_dat_o[23] = net178;
 assign wbs_dat_o[24] = net179;
 assign wbs_dat_o[25] = net180;
 assign wbs_dat_o[26] = net181;
 assign wbs_dat_o[27] = net182;
 assign wbs_dat_o[28] = net183;
 assign wbs_dat_o[29] = net184;
 assign wbs_dat_o[2] = net157;
 assign wbs_dat_o[30] = net185;
 assign wbs_dat_o[31] = net186;
 assign wbs_dat_o[3] = net158;
 assign wbs_dat_o[4] = net159;
 assign wbs_dat_o[5] = net160;
 assign wbs_dat_o[6] = net161;
 assign wbs_dat_o[7] = net162;
 assign wbs_dat_o[8] = net163;
 assign wbs_dat_o[9] = net164;
endmodule
